package encoderr;
class transaction;
rand bit rst;
rand bit [3:0] D;
function new();
endfunction
endclass
endpackage

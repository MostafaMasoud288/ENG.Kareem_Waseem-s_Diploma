package shared_pck;

typedef enum  {SHIFT,ROTATE} mode_e;

typedef enum  {RIGHT,LEFT} direction_e;

endpackage
